VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.5 ;
  WIDTH 0.2 ;
END M1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.5 ;
  WIDTH 0.2 ;
END M2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.5 ;
  WIDTH 0.2 ;
END M3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.5 ;
  WIDTH 0.2 ;
END M4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.5 ;
  WIDTH 0.2 ;
END M5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.5 ;
  WIDTH 0.2 ;
END M6

MACRO NAND2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.0 BY 4.0 ;
  SYMMETRY X Y ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.4 1.0 0.6 1.2 ;  # Center 0.5 (Aligned!)
    END
  END
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.4 2.0 0.6 2.2 ;  # Center 0.5 (Aligned!)
    END
  END
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 1.4 2.0 1.6 2.2 ;  # Center 1.5 (Aligned!)
    END
  END
END NAND2

MACRO DFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.0 BY 4.0 ;
  SYMMETRY X Y ;
  SITE CORE ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.4 1.0 0.6 1.2 ;
    END
  END
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT 3.4 1.0 3.6 1.2 ;
    END
  END
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT 0.4 3.0 0.6 3.2 ;
    END
  END
END DFF

END LIBRARY
